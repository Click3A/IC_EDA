interface intf(input logic clk,reset);
    logic [3:0]a;
    logic [3:0]b;
    logic [7:0]c;
endinterface
