class generator;
    rand transaction trans;

    mailbox gen2driv;

    int repeat_time;

    function new(mailbox gen2driv);
        this.gen2driv = gen2driv;
    endfunction

    task main();
        repeat(repeat_time)begin
            trans = new();
            trans.randomize();
            gen2driv.put(trans);
        end
    endtask
endclass
